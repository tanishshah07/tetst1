`include "mux.v"
module top;
wire out;
reg [1:0] i;
reg s;
mux dut(out,i,s);
initial begin
	repeat(5) begin
		#7
	{i,s}=$random;
	$display("out=%b,i=%b,s=%b",out,i,s);
end
end
endmodule
